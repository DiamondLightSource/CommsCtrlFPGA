----------------------------------------------------------------------
--  Project      : Diamond FOFB Communication Controller
--  Filename     :
--  Purpose      : Virtex2Pro MGT interface
--  Responsible  : Isa S. Uzun
----------------------------------------------------------------------
--  Copyright (c) 2007 Diamond Light Source Ltd.
--  All rights reserved.
----------------------------------------------------------------------
--  Description: This is the top-level interface module that instantiates
--  MGT Tile and user logic to interface CC.
----------------------------------------------------------------------
--  Limitations & Assumptions:
----------------------------------------------------------------------
--  Known Errors: Please send any bug reports to isa.uzun@diamond.ac.uk
----------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

library work;
use work.fofb_cc_pkg.all;

entity fofb_cc_mgt_if is
    generic (
        -- CC Design selection parameters
        DEVICE                  : device_t := BPM;
        LaneCount               : integer := 4;
        TX_IDLE_NUM             : natural := 16;    --32767 cc
        RX_IDLE_NUM             : natural := 13;    --4095 cc
        SEND_ID_NUM             : natural := 14     --8191 cc
    );
    port (
        -- clocks and resets
        refclk_i                : in  std_logic;
        userclk_i               : in  std_logic;
        mgtreset_i              : in  std_logic;

        rxn_i                   : in  std_logic_vector(LaneCount-1 downto 0);
        rxp_i                   : in  std_logic_vector(LaneCount-1 downto 0);
        txn_o                   : out std_logic_vector(LaneCount-1 downto 0);
        txp_o                   : out std_logic_vector(LaneCount-1 downto 0);

        -- time frame sync
        timeframe_start_i       : in  std_logic;
        timeframe_end_i         : in  std_logic;
        timeframe_val_i         : in  std_logic_vector(15 downto 0);
        bpmid_i                 : in  std_logic_vector(7 downto 0);

        -- mgt configuration 
        powerdown_i             : in  std_logic_vector(3 downto 0);
        loopback_i              : in  std_logic_vector(7 downto 0);

        -- status information
        linksup_o               : out std_logic_vector(7 downto 0);
        frameerror_cnt_o        : inout std_logic_2d_16(3 downto 0); 
        softerror_cnt_o         : inout std_logic_2d_16(3 downto 0); 
        harderror_cnt_o         : inout std_logic_2d_16(3 downto 0); 
        txpck_cnt_o             : out std_logic_2d_16(3 downto 0);
        rxpck_cnt_o             : out std_logic_2d_16(3 downto 0);

        -- network information
        tfs_bit_o               : out std_logic_vector(3 downto 0);
        link_partner_o          : out std_logic_2d_10(3 downto 0);
        pmc_timeframe_val_o     : out std_logic_2d_16(3 downto 0);
        pmc_timestamp_val_o     : out std_logic_2d_32(3 downto 0);

        -- tx/rx state machine status for reset operation
        tx_sm_busy_o            : out std_logic_vector(LaneCount-1 downto 0);
        rx_sm_busy_o            : out std_logic_vector(LaneCount-1 downto 0);

        -- TX FIFO interface
        tx_dat_i                : in  std_logic_2d_16(LaneCount-1 downto 0);
        txf_empty_i             : in  std_logic_vector(LaneCount-1 downto 0);
        txf_rd_en_o             : out std_logic_vector(LaneCount-1 downto 0);

        -- RX FIFO interface
        rxf_full_i              : in  std_logic_vector(LaneCount-1 downto 0);
        rx_dat_o                : out std_logic_2d_16(LaneCount-1 downto 0);
        rx_dat_val_o            : out std_logic_vector(LaneCount-1 downto 0)
    );
end fofb_cc_mgt_if;

architecture rtl of fofb_cc_mgt_if is 

signal txdata               : std_logic_2d_16(LaneCount-1 downto 0);
signal rxdata               : std_logic_2d_16(LaneCount-1 downto 0);
signal txcharisk            : std_logic_2d_2(LaneCount-1 downto 0);
signal rxcharisk            : std_logic_2d_2(LaneCount-1 downto 0);
signal encommaalign         : std_logic_vector(LaneCount-1 downto 0);
signal txkerr               : std_logic_2d_2(LaneCount-1 downto 0);
signal txbuferr             : std_logic_vector(LaneCount-1 downto 0);
signal rxbuferr             : std_logic_vector(LaneCount-1 downto 0);
signal rxrealign            : std_logic_vector(LaneCount-1 downto 0);
signal rxdisperr            : std_logic_2d_2(LaneCount-1 downto 0);
signal rxnotintable         : std_logic_2d_2(LaneCount-1 downto 0);
signal rxreset              : std_logic_vector(LaneCount-1 downto 0);
signal txreset              : std_logic_vector(LaneCount-1 downto 0);
signal rxcheckingcrc        : std_logic_vector(LaneCount-1 downto 0);
signal rxcrcerr             : std_logic_vector(LaneCount-1 downto 0);
signal refclksel            : std_logic;

begin

refclksel <= '0'; -- for BREFCLK

MGT_IF_GEN: for N in 0 to (LaneCount-1) generate

MGT_LANES: entity work.fofb_cc_mgt_lane
    generic map(
        -- CC Design selection parameters
        TX_IDLE_NUM             => TX_IDLE_NUM,
        RX_IDLE_NUM             => RX_IDLE_NUM,
        SEND_ID_NUM             => SEND_ID_NUM
    )
    port map (
        userclk_i               => userclk_i,
        mgtreset_i              => mgtreset_i,
        rxreset_o               => rxreset(N),
        txreset_o               => txreset(N),
        powerdown_i             => powerdown_i(N),

        timeframe_start_i       => timeframe_start_i,
        timeframe_end_i         => timeframe_end_i,
        timeframe_val_i         => timeframe_val_i,
        bpmid_i                 => bpmid_i,

        linksup_o               => linksup_o(2*N+1 downto 2*N),
        frameerror_cnt_o        => frameerror_cnt_o(N),
        softerror_cnt_o         => softerror_cnt_o(N),
        harderror_cnt_o         => harderror_cnt_o(N),
        txpck_cnt_o             => txpck_cnt_o(N),
        rxpck_cnt_o             => rxpck_cnt_o(N),

        tfs_bit_o               => tfs_bit_o(N),
        link_partner_o          => link_partner_o(N),
        pmc_timeframe_val_o     => pmc_timeframe_val_o(N),
        timestamp_val_o         => pmc_timestamp_val_o(N),

        tx_sm_busy_o            => tx_sm_busy_o(N),
        rx_sm_busy_o            => rx_sm_busy_o(N),

        tx_dat_i                => tx_dat_i(N),
        txf_empty_i             => txf_empty_i(N),
        txf_rd_en_o             => txf_rd_en_o(N),

        rxf_full_i              => rxf_full_i(N),
        rx_dat_o                => rx_dat_o(N),
        rx_dat_val_o            => rx_dat_val_o(N),

        txdata_o                => txdata(N),
        txcharisk_o             => txcharisk(N),
        rxdata_i                => rxdata(N),
        rxcharisk_i             => rxcharisk(N),
        encommaalign_o          => encommaalign(N),
        txkerr_i                => txkerr(N),
        txbuferr_i              => txbuferr(N),
        rxbuferr_i              => rxbuferr(N),
        rxrealign_i             => rxrealign(N),
        rxdisperr_i             => rxdisperr(N),
        rxnotintable_i          => rxnotintable(N),
        rxcrcerr_i              => rxcrcerr(N),
        rxcheckingcrc_i         => rxcheckingcrc(N)
    );

MGT_TILES : entity work.fofb_cc_mgt_tile
    port map (
        brefclk_i               => refclk_i,
        refclksel_i             => refclksel,
        userclk_i               => userclk_i,
        encommaalign_i          => encommaalign(N),
        loopback_i              => loopback_i(2*N+1 downto 2*N),
        powerdown_i             => powerdown_i(N),
        rxn_i                   => rxn_i(N),
        rxp_i                   => rxp_i(N),
        rxreset_i               => rxreset(N),
        txcharisk_i             => txcharisk(N),
        txdata_i                => txdata(N),
        txreset_i               => txreset(N),
        rxbufstatus_o           => rxbuferr(N),
        rxcharisk_o             => rxcharisk(N),
        rxcheckingcrc_o         => rxcheckingcrc(N),
        rxcrcerr_o              => rxcrcerr(N),
        rxdata_o                => rxdata(N),
        rxdisperr_o             => rxdisperr(N),
        rxnotintable_o          => rxnotintable(N),
        rxrealign_o             => rxrealign(N),
        txbuferr_o              => txbuferr(N),
        txkerr_o                => txkerr(N),
        txn_o                   => txn_o(N),
        txp_o                   => txp_o(N)
);

end generate;

end rtl;
