library ieee;
use ieee.std_logic_1164.all;
package fofb_cc_version is
constant FPGAFirmwareVersion: std_logic_vector(31 downto 0) := X"00003004";
end fofb_cc_version;
