entity cdc_ctrl is
end;

architecture ctrl of cdc_ctrl is
begin

-- 0in set_cdc_clock refclk_p_i -period 8
-- 0in set_cdc_clock refclk_n_i -period 8
-- 0in set_cdc_clock adcclk_i   -period 8
-- 0in set_cdc_clock sysclk_i   -period 8

end ctrl;

