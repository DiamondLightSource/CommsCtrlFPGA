-------------------------------------------------------------------------------
--$Date: 2008/04/01 22:44:07 $
--$RCSfile: sim_reset_mgt_model_vhd.ejava,v $
--$Revision: 1.1.2.2 $
--------------------------------------------------------------------------------
--   ____  ____ 
--  /   /\/   / 
-- /___/  \  /    Vendor: Xilinx 
-- \   \   \/     Version : 1.9
--  \   \         Application : GTP Wizard
--  /   /         Filename : sim_reset_mgt_model.vhd
-- /___/   /\     Timestamp : 
-- \   \  /  \ 
--  \___\/\___\ 
--
--
-- Module SIM_RESET_MGT_MODEL
-- Generated by Xilinx RocketIO Wizard
--
-- The Reset On Configuration(ROC) module is part of the UNISIM library
-- and is required for emulating the GSR pulse at the beginning of functional
-- simulation in order to correctly reset the VHDL MGT smart model.This module
-- is required for simulation only.


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library UNISIM;
use UNISIM.VCOMPONENTS.ALL;

--***************************** Entity Declaration *****************************

entity SIM_RESET_MGT_MODEL is
port 
(
    GSR_IN     : in std_logic
);
end SIM_RESET_MGT_MODEL;

architecture BEHAVIORAL of SIM_RESET_MGT_MODEL is
  
                  
--********************************* Main Body of Code****************************
                       
begin                      
    GSR <= GSR_IN;                       
    ------------------------------  ROCBUF Instantiation -----------------------   
    -- This component is required for correctly resetting the VHDL GTP component on configuration
    -- It is for simulation alone and will be ripped out during synthesis.
    U1 : ROCBUF 
    port map 
    (
        I => GSR,
        O => open
    ); 


end BEHAVIORAL;

